// Benchmark "top" written by ABC on Tue Apr 15 22:49:29 2025

module top ( 
    pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9, pi10,
    po0, po1, po2, po3, po4  );
  input  pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9, pi10;
  output po0, po1, po2, po3, po4;
  wire new_new_n16, new_new_n15, new_new_n17, new_new_n14, new_new_n18,
    new_new_n13, new_new_n19, new_new_n11, new_new_n12, new_new_n20,
    new_new_n25, new_new_n24, new_new_n26, new_new_n23, new_new_n27,
    new_new_n22, new_new_n28, new_new_n21, new_new_n29, new_new_n37,
    new_new_n36, new_new_n38, new_new_n34, new_new_n35, new_new_n39,
    new_new_n32, new_new_n33, new_new_n40, new_new_n30, new_new_n31,
    new_new_n41, new_new_n46, new_new_n45, new_new_n47, new_new_n44,
    new_new_n48, new_new_n43, new_new_n49, new_new_n42, new_new_n50,
    new_new_n55, new_new_n54, new_new_n56, new_new_n53, new_new_n57,
    new_new_n52, new_new_n58, new_new_n51, new_new_n59;
  assign new_new_n16 = pi1 & pi6;
  assign new_new_n15 = pi5 & pi7;
  assign new_new_n17 = ~new_new_n16 ^ ~new_new_n15;
  assign new_new_n14 = pi4 & pi8;
  assign new_new_n18 = ~new_new_n17 ^ ~new_new_n14;
  assign new_new_n13 = pi3 & pi9;
  assign new_new_n19 = ~new_new_n18 ^ ~new_new_n13;
  assign new_new_n11 = ~pi5 ^ ~pi2;
  assign new_new_n12 = pi10 & new_new_n11;
  assign new_new_n20 = ~new_new_n19 ^ ~new_new_n12;
  assign new_new_n25 = pi2 & pi6;
  assign new_new_n24 = pi1 & pi7;
  assign new_new_n26 = ~new_new_n25 ^ ~new_new_n24;
  assign new_new_n23 = pi5 & pi8;
  assign new_new_n27 = ~new_new_n26 ^ ~new_new_n23;
  assign new_new_n22 = pi4 & pi9;
  assign new_new_n28 = ~new_new_n27 ^ ~new_new_n22;
  assign new_new_n21 = pi3 & pi10;
  assign new_new_n29 = ~new_new_n28 ^ ~new_new_n21;
  assign new_new_n37 = pi3 & pi6;
  assign new_new_n36 = pi7 & new_new_n11;
  assign new_new_n38 = ~new_new_n37 ^ ~new_new_n36;
  assign new_new_n34 = ~pi4 ^ ~pi1;
  assign new_new_n35 = pi8 & new_new_n34;
  assign new_new_n39 = ~new_new_n38 ^ ~new_new_n35;
  assign new_new_n32 = ~pi5 ^ ~pi3;
  assign new_new_n33 = pi9 & new_new_n32;
  assign new_new_n40 = ~new_new_n39 ^ ~new_new_n33;
  assign new_new_n30 = ~new_new_n11 ^ ~pi4;
  assign new_new_n31 = pi10 & new_new_n30;
  assign new_new_n41 = ~new_new_n40 ^ ~new_new_n31;
  assign new_new_n46 = pi4 & pi6;
  assign new_new_n45 = pi3 & pi7;
  assign new_new_n47 = ~new_new_n46 ^ ~new_new_n45;
  assign new_new_n44 = pi8 & new_new_n11;
  assign new_new_n48 = ~new_new_n47 ^ ~new_new_n44;
  assign new_new_n43 = pi9 & new_new_n34;
  assign new_new_n49 = ~new_new_n48 ^ ~new_new_n43;
  assign new_new_n42 = pi10 & new_new_n32;
  assign new_new_n50 = ~new_new_n49 ^ ~new_new_n42;
  assign new_new_n55 = pi5 & pi6;
  assign new_new_n54 = pi4 & pi7;
  assign new_new_n56 = ~new_new_n55 ^ ~new_new_n54;
  assign new_new_n53 = pi3 & pi8;
  assign new_new_n57 = ~new_new_n56 ^ ~new_new_n53;
  assign new_new_n52 = pi9 & new_new_n11;
  assign new_new_n58 = ~new_new_n57 ^ ~new_new_n52;
  assign new_new_n51 = pi10 & new_new_n34;
  assign new_new_n59 = ~new_new_n58 ^ ~new_new_n51;
  assign po0 = new_new_n20;
  assign po1 = new_new_n29;
  assign po2 = new_new_n41;
  assign po3 = new_new_n50;
  assign po4 = new_new_n59;
endmodule


